module Compute_S
(
  input  wire [(`N*`SYMBOL_WIDTH)-1:0] v,
  output wire [`SYMBOL_WIDTH-1:0]      s1,
  output wire [`SYMBOL_WIDTH-1:0]      s2
);
  
  wire  [143:0] H_row_0;
  wire  [143:0] H_row_1;
  wire  [143:0] H_row_2;
  wire  [143:0] H_row_3;
  wire  [143:0] H_row_4;
  wire  [143:0] H_row_5;
  wire  [143:0] H_row_6;
  wire  [143:0] H_row_7;
  wire  [143:0] H_row_8;
  wire  [143:0] H_row_9;
  wire  [143:0] H_row_10;
  wire  [143:0] H_row_11;
  wire  [143:0] H_row_12;
  wire  [143:0] H_row_13;
  wire  [143:0] H_row_14;
  wire  [143:0] H_row_15;
           
      assign H_row_0  = 144'b000100000000110000000111111001111101110010001111100110111110110000101100101110001100111100011111100001111111011111000000100001001000000000000000;
      assign H_row_1  = 144'b000010000000011010111011110010110110111011111111111101010111011000010110010111001101111110110111111110111100001101100000010000100100000000000000;
      assign H_row_2  = 144'b000001000000001111100101110111010011011111000111110000100011101100001011001011101101011111100011110001011101100100110000001000010010000000000000;
      assign H_row_3  = 144'b000000101011100111001010110101101010001111011011011000011010010110111101000101111101001111001001110110101101010000011000101010000001000000000000;
      assign H_row_4  = 144'b000000011110010001100101011010111110100111010101100010001110101011100110101100111101000111011100011011010110101000001100010101000000100000000000;
      assign H_row_5  = 144'b101110000111001010001010100011011100110011010010010001000111010101110011111000011101000001101110100011100011010100000110001010100000010000000000;
      assign H_row_6  = 144'b010111000011100101000101111111100110011001101001001000101000001010000001110010000110100000110111010001111010001000000011000101010000001000000000;
      assign H_row_7  = 144'b001011101010010010011010011111110011001110001100000100010100000111111000011001000011010010100011100110110101000110111001101100100000000100000000;
      assign H_row_8  = 144'b011000000011100000011110101101111100110101101101010001100001000100000100001011111111100010001101100111100101011110010101010010110000000010000000;
      assign H_row_9  = 144'b001100000001110000001111111000111101111010001110001000111011000000000010101011110111110011111110010011111001001111110010100111010000000001000000;
      assign H_row_10 = 144'b000110000000111010111111110010010110111101000111101010010101100000000001111011110011111001111111100111111111000101111001111101100000000000100000;
      assign H_row_11 = 144'b000011000000011111100111110111001000111110011011111011000010110010111000110011110001111110000111111101111100000010000100011110110000000000010000;
      assign H_row_12 = 144'b000001101011101111001011011011101111111111110101011101100001011001011100110111111011011111111011110000110110000001000010100001010000000000001000;
      assign H_row_13 = 144'b000000111110010111011101001101111100011111000010001110110000101100101110110101111110001111000101110110010011000000100001111110100000000000000100;
      assign H_row_14 = 144'b101110011100101011010110101000111101101101100001101001011011110100010111110100111100100111011010110101000001100010101000011111010000000000000010;
      assign H_row_15 = 144'b111001000110010101101011111010011101010110001000111010101110011010110011110100011101110001101101011010100000110001010100100001100000000000000001;
      
  assign s1[0] = ^(v & H_row_0)  ;
  assign s1[1] = ^(v & H_row_1)  ;
  assign s1[2] = ^(v & H_row_2)  ;
  assign s1[3] = ^(v & H_row_3)  ;
  assign s1[4] = ^(v & H_row_4)  ;
  assign s1[5] = ^(v & H_row_5)  ;
  assign s1[6] = ^(v & H_row_6)  ;
  assign s1[7] = ^(v & H_row_7)  ;
  assign s2[0] = ^(v & H_row_8)  ;
  assign s2[1] = ^(v & H_row_9)  ;
  assign s2[2] = ^(v & H_row_10) ;
  assign s2[3] = ^(v & H_row_11) ;
  assign s2[4] = ^(v & H_row_12) ;
  assign s2[5] = ^(v & H_row_13) ;
  assign s2[6] = ^(v & H_row_14) ;
  assign s2[7] = ^(v & H_row_15) ;
  
endmodule
