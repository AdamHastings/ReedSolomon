module Compute_S
(
  input  wire [(`N*`SYMBOL_WIDTH)-1:0] v,
  output wire [`SYMBOL_WIDTH-1:0]      s1,
  output wire [`SYMBOL_WIDTH-1:0]      s2
);
  
  wire  [143:0] H_row_0;
  wire  [143:0] H_row_1;
  wire  [143:0] H_row_2;
  wire  [143:0] H_row_3;
  wire  [143:0] H_row_4;
  wire  [143:0] H_row_5;
           
      assign H_row_0  = 144'b000100000000110000000111111001111101110010001111100110111110110000101100101110001100111100011111100001111111011111000000100001001000000000000000;
      assign H_row_1  = 144'b000010000000011010111011110010110110111011111111111101010111011000010110010111001101111110110111111110111100001101100000010000100100000000000000;
      assign H_row_2  = 144'b000001000000001111100101110111010011011111000111110000100011101100001011001011101101011111100011110001011101100100110000001000010010000000000000;
      assign H_row_3  = 144'b000000101011100111001010110101101010001111011011011000011010010110111101000101111101001111001001110110101101010000011000101010000001000000000000;
      assign H_row_4  = 144'b000000011110010001100101011010111110100111010101100010001110101011100110101100111101000111011100011011010110101000001100010101000000100000000000;
      assign H_row_5  = 144'b101110000111001010001010100011011100110011010010010001000111010101110011111000011101000001101110100011100011010100000110001010100000010000000000;
      
  assign s1[0] = ^(v & H_row_0)  ;
  assign s1[1] = ^(v & H_row_1)  ;
  assign s1[2] = ^(v & H_row_2)  ;
  assign s2[0] = ^(v & H_row_8)  ;
  assign s2[1] = ^(v & H_row_9)  ;
  assign s2[2] = ^(v & H_row_10) ;
  
endmodule
