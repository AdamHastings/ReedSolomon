`define SYMBOL_WIDTH 8
`define N 18
`define K 16

module Symbol_Lookup
(
  input   wire [`SYMBOL_WIDTH-1:0] in,
  output  reg  [`SYMBOL_WIDTH-1:0] out
);
  always @* begin
    case(in)
      8'd0 : out <= 8'b00000000;
      8'd1 : out <= 8'b10000000;
      8'd2 : out <= 8'b01000000;
      8'd3 : out <= 8'b00100000;
      8'd4 : out <= 8'b00010000;
      8'd5 : out <= 8'b00001000;
      8'd6 : out <= 8'b00000100;
      8'd7 : out <= 8'b00000010;
      8'd8 : out <= 8'b00000001;
      8'd9 : out <= 8'b10111000;
      8'd10 : out <= 8'b01011100;
      8'd11 : out <= 8'b00101110;
      8'd12 : out <= 8'b00010111;
      8'd13 : out <= 8'b10110011;
      8'd14 : out <= 8'b11100001;
      8'd15 : out <= 8'b11001000;
      8'd16 : out <= 8'b01100100;
      8'd17 : out <= 8'b00110010;
      8'd18 : out <= 8'b00011001;
      8'd19 : out <= 8'b10110100;
      8'd20 : out <= 8'b01011010;
      8'd21 : out <= 8'b00101101;
      8'd22 : out <= 8'b10101110;
      8'd23 : out <= 8'b01010111;
      8'd24 : out <= 8'b10010011;
      8'd25 : out <= 8'b11110001;
      8'd26 : out <= 8'b11000000;
      8'd27 : out <= 8'b01100000;
      8'd28 : out <= 8'b00110000;
      8'd29 : out <= 8'b00011000;
      8'd30 : out <= 8'b00001100;
      8'd31 : out <= 8'b00000110;
      8'd32 : out <= 8'b00000011;
      8'd33 : out <= 8'b10111001;
      8'd34 : out <= 8'b11100100;
      8'd35 : out <= 8'b01110010;
      8'd36 : out <= 8'b00111001;
      8'd37 : out <= 8'b10100100;
      8'd38 : out <= 8'b01010010;
      8'd39 : out <= 8'b00101001;
      8'd40 : out <= 8'b10101100;
      8'd41 : out <= 8'b01010110;
      8'd42 : out <= 8'b00101011;
      8'd43 : out <= 8'b10101101;
      8'd44 : out <= 8'b11101110;
      8'd45 : out <= 8'b01110111;
      8'd46 : out <= 8'b10000011;
      8'd47 : out <= 8'b11111001;
      8'd48 : out <= 8'b11000100;
      8'd49 : out <= 8'b01100010;
      8'd50 : out <= 8'b00110001;
      8'd51 : out <= 8'b10100000;
      8'd52 : out <= 8'b01010000;
      8'd53 : out <= 8'b00101000;
      8'd54 : out <= 8'b00010100;
      8'd55 : out <= 8'b00001010;
      8'd56 : out <= 8'b00000101;
      8'd57 : out <= 8'b10111010;
      8'd58 : out <= 8'b01011101;
      8'd59 : out <= 8'b10010110;
      8'd60 : out <= 8'b01001011;
      8'd61 : out <= 8'b10011101;
      8'd62 : out <= 8'b11110110;
      8'd63 : out <= 8'b01111011;
      8'd64 : out <= 8'b10000101;
      8'd65 : out <= 8'b11111010;
      8'd66 : out <= 8'b01111101;
      8'd67 : out <= 8'b10000110;
      8'd68 : out <= 8'b01000011;
      8'd69 : out <= 8'b10011001;
      8'd70 : out <= 8'b11110100;
      8'd71 : out <= 8'b01111010;
      8'd72 : out <= 8'b00111101;
      8'd73 : out <= 8'b10100110;
      8'd74 : out <= 8'b01010011;
      8'd75 : out <= 8'b10010001;
      8'd76 : out <= 8'b11110000;
      8'd77 : out <= 8'b01111000;
      8'd78 : out <= 8'b00111100;
      8'd79 : out <= 8'b00011110;
      8'd80 : out <= 8'b00001111;
      8'd81 : out <= 8'b10111111;
      8'd82 : out <= 8'b11100111;
      8'd83 : out <= 8'b11001011;
      8'd84 : out <= 8'b11011101;
      8'd85 : out <= 8'b11010110;
      8'd86 : out <= 8'b01101011;
      8'd87 : out <= 8'b10001101;
      8'd88 : out <= 8'b11111110;
      8'd89 : out <= 8'b01111111;
      8'd90 : out <= 8'b10000111;
      8'd91 : out <= 8'b11111011;
      8'd92 : out <= 8'b11000101;
      8'd93 : out <= 8'b11011010;
      8'd94 : out <= 8'b01101101;
      8'd95 : out <= 8'b10001110;
      8'd96 : out <= 8'b01000111;
      8'd97 : out <= 8'b10011011;
      8'd98 : out <= 8'b11110101;
      8'd99 : out <= 8'b11000010;
      8'd100 : out <= 8'b01100001;
      8'd101 : out <= 8'b10001000;
      8'd102 : out <= 8'b01000100;
      8'd103 : out <= 8'b00100010;
      8'd104 : out <= 8'b00010001;
      8'd105 : out <= 8'b10110000;
      8'd106 : out <= 8'b01011000;
      8'd107 : out <= 8'b00101100;
      8'd108 : out <= 8'b00010110;
      8'd109 : out <= 8'b00001011;
      8'd110 : out <= 8'b10111101;
      8'd111 : out <= 8'b11100110;
      8'd112 : out <= 8'b01110011;
      8'd113 : out <= 8'b10000001;
      8'd114 : out <= 8'b11111000;
      8'd115 : out <= 8'b01111100;
      8'd116 : out <= 8'b00111110;
      8'd117 : out <= 8'b00011111;
      8'd118 : out <= 8'b10110111;
      8'd119 : out <= 8'b11100011;
      8'd120 : out <= 8'b11001001;
      8'd121 : out <= 8'b11011100;
      8'd122 : out <= 8'b01101110;
      8'd123 : out <= 8'b00110111;
      8'd124 : out <= 8'b10100011;
      8'd125 : out <= 8'b11101001;
      8'd126 : out <= 8'b11001100;
      8'd127 : out <= 8'b01100110;
      8'd128 : out <= 8'b00110011;
      8'd129 : out <= 8'b10100001;
      8'd130 : out <= 8'b11101000;
      8'd131 : out <= 8'b01110100;
      8'd132 : out <= 8'b00111010;
      8'd133 : out <= 8'b00011101;
      8'd134 : out <= 8'b10110110;
      8'd135 : out <= 8'b01011011;
      8'd136 : out <= 8'b10010101;
      8'd137 : out <= 8'b11110010;
      8'd138 : out <= 8'b01111001;
      8'd139 : out <= 8'b10000100;
      8'd140 : out <= 8'b01000010;
      8'd141 : out <= 8'b00100001;
      8'd142 : out <= 8'b10101000;
      8'd143 : out <= 8'b01010100;
      8'd144 : out <= 8'b00101010;
      8'd145 : out <= 8'b00010101;
      8'd146 : out <= 8'b10110010;
      8'd147 : out <= 8'b01011001;
      8'd148 : out <= 8'b10010100;
      8'd149 : out <= 8'b01001010;
      8'd150 : out <= 8'b00100101;
      8'd151 : out <= 8'b10101010;
      8'd152 : out <= 8'b01010101;
      8'd153 : out <= 8'b10010010;
      8'd154 : out <= 8'b01001001;
      8'd155 : out <= 8'b10011100;
      8'd156 : out <= 8'b01001110;
      8'd157 : out <= 8'b00100111;
      8'd158 : out <= 8'b10101011;
      8'd159 : out <= 8'b11101101;
      8'd160 : out <= 8'b11001110;
      8'd161 : out <= 8'b01100111;
      8'd162 : out <= 8'b10001011;
      8'd163 : out <= 8'b11111101;
      8'd164 : out <= 8'b11000110;
      8'd165 : out <= 8'b01100011;
      8'd166 : out <= 8'b10001001;
      8'd167 : out <= 8'b11111100;
      8'd168 : out <= 8'b01111110;
      8'd169 : out <= 8'b00111111;
      8'd170 : out <= 8'b10100111;
      8'd171 : out <= 8'b11101011;
      8'd172 : out <= 8'b11001101;
      8'd173 : out <= 8'b11011110;
      8'd174 : out <= 8'b01101111;
      8'd175 : out <= 8'b10001111;
      8'd176 : out <= 8'b11111111;
      8'd177 : out <= 8'b11000111;
      8'd178 : out <= 8'b11011011;
      8'd179 : out <= 8'b11010101;
      8'd180 : out <= 8'b11010010;
      8'd181 : out <= 8'b01101001;
      8'd182 : out <= 8'b10001100;
      8'd183 : out <= 8'b01000110;
      8'd184 : out <= 8'b00100011;
      8'd185 : out <= 8'b10101001;
      8'd186 : out <= 8'b11101100;
      8'd187 : out <= 8'b01110110;
      8'd188 : out <= 8'b00111011;
      8'd189 : out <= 8'b10100101;
      8'd190 : out <= 8'b11101010;
      8'd191 : out <= 8'b01110101;
      8'd192 : out <= 8'b10000010;
      8'd193 : out <= 8'b01000001;
      8'd194 : out <= 8'b10011000;
      8'd195 : out <= 8'b01001100;
      8'd196 : out <= 8'b00100110;
      8'd197 : out <= 8'b00010011;
      8'd198 : out <= 8'b10110001;
      8'd199 : out <= 8'b11100000;
      8'd200 : out <= 8'b01110000;
      8'd201 : out <= 8'b00111000;
      8'd202 : out <= 8'b00011100;
      8'd203 : out <= 8'b00001110;
      8'd204 : out <= 8'b00000111;
      8'd205 : out <= 8'b10111011;
      8'd206 : out <= 8'b11100101;
      8'd207 : out <= 8'b11001010;
      8'd208 : out <= 8'b01100101;
      8'd209 : out <= 8'b10001010;
      8'd210 : out <= 8'b01000101;
      8'd211 : out <= 8'b10011010;
      8'd212 : out <= 8'b01001101;
      8'd213 : out <= 8'b10011110;
      8'd214 : out <= 8'b01001111;
      8'd215 : out <= 8'b10011111;
      8'd216 : out <= 8'b11110111;
      8'd217 : out <= 8'b11000011;
      8'd218 : out <= 8'b11011001;
      8'd219 : out <= 8'b11010100;
      8'd220 : out <= 8'b01101010;
      8'd221 : out <= 8'b00110101;
      8'd222 : out <= 8'b10100010;
      8'd223 : out <= 8'b01010001;
      8'd224 : out <= 8'b10010000;
      8'd225 : out <= 8'b01001000;
      8'd226 : out <= 8'b00100100;
      8'd227 : out <= 8'b00010010;
      8'd228 : out <= 8'b00001001;
      8'd229 : out <= 8'b10111100;
      8'd230 : out <= 8'b01011110;
      8'd231 : out <= 8'b00101111;
      8'd232 : out <= 8'b10101111;
      8'd233 : out <= 8'b11101111;
      8'd234 : out <= 8'b11001111;
      8'd235 : out <= 8'b11011111;
      8'd236 : out <= 8'b11010111;
      8'd237 : out <= 8'b11010011;
      8'd238 : out <= 8'b11010001;
      8'd239 : out <= 8'b11010000;
      8'd240 : out <= 8'b01101000;
      8'd241 : out <= 8'b00110100;
      8'd242 : out <= 8'b00011010;
      8'd243 : out <= 8'b00001101;
      8'd244 : out <= 8'b10111110;
      8'd245 : out <= 8'b01011111;
      8'd246 : out <= 8'b10010111;
      8'd247 : out <= 8'b11110011;
      8'd248 : out <= 8'b11000001;
      8'd249 : out <= 8'b11011000;
      8'd250 : out <= 8'b01101100;
      8'd251 : out <= 8'b00110110;
      8'd252 : out <= 8'b00011011;
      8'd253 : out <= 8'b10110101;
      8'd254 : out <= 8'b11100010;
      8'd255 : out <= 8'b01110001;
      default: out <= 8'b00000000;
    endcase
  end
endmodule

module Index_Lookup
(
  input   wire [`SYMBOL_WIDTH-1:0] in,
  output  reg  [`SYMBOL_WIDTH-1:0] out
);
  always @* begin
    case(in)
      8'b00000000 : out <= 8'd0;
      8'b10000000 : out <= 8'd1;
      8'b01000000 : out <= 8'd2;
      8'b00100000 : out <= 8'd3;
      8'b00010000 : out <= 8'd4;
      8'b00001000 : out <= 8'd5;
      8'b00000100 : out <= 8'd6;
      8'b00000010 : out <= 8'd7;
      8'b00000001 : out <= 8'd8;
      8'b10111000 : out <= 8'd9;
      8'b01011100 : out <= 8'd10;
      8'b00101110 : out <= 8'd11;
      8'b00010111 : out <= 8'd12;
      8'b10110011 : out <= 8'd13;
      8'b11100001 : out <= 8'd14;
      8'b11001000 : out <= 8'd15;
      8'b01100100 : out <= 8'd16;
      8'b00110010 : out <= 8'd17;
      8'b00011001 : out <= 8'd18;
      8'b10110100 : out <= 8'd19;
      8'b01011010 : out <= 8'd20;
      8'b00101101 : out <= 8'd21;
      8'b10101110 : out <= 8'd22;
      8'b01010111 : out <= 8'd23;
      8'b10010011 : out <= 8'd24;
      8'b11110001 : out <= 8'd25;
      8'b11000000 : out <= 8'd26;
      8'b01100000 : out <= 8'd27;
      8'b00110000 : out <= 8'd28;
      8'b00011000 : out <= 8'd29;
      8'b00001100 : out <= 8'd30;
      8'b00000110 : out <= 8'd31;
      8'b00000011 : out <= 8'd32;
      8'b10111001 : out <= 8'd33;
      8'b11100100 : out <= 8'd34;
      8'b01110010 : out <= 8'd35;
      8'b00111001 : out <= 8'd36;
      8'b10100100 : out <= 8'd37;
      8'b01010010 : out <= 8'd38;
      8'b00101001 : out <= 8'd39;
      8'b10101100 : out <= 8'd40;
      8'b01010110 : out <= 8'd41;
      8'b00101011 : out <= 8'd42;
      8'b10101101 : out <= 8'd43;
      8'b11101110 : out <= 8'd44;
      8'b01110111 : out <= 8'd45;
      8'b10000011 : out <= 8'd46;
      8'b11111001 : out <= 8'd47;
      8'b11000100 : out <= 8'd48;
      8'b01100010 : out <= 8'd49;
      8'b00110001 : out <= 8'd50;
      8'b10100000 : out <= 8'd51;
      8'b01010000 : out <= 8'd52;
      8'b00101000 : out <= 8'd53;
      8'b00010100 : out <= 8'd54;
      8'b00001010 : out <= 8'd55;
      8'b00000101 : out <= 8'd56;
      8'b10111010 : out <= 8'd57;
      8'b01011101 : out <= 8'd58;
      8'b10010110 : out <= 8'd59;
      8'b01001011 : out <= 8'd60;
      8'b10011101 : out <= 8'd61;
      8'b11110110 : out <= 8'd62;
      8'b01111011 : out <= 8'd63;
      8'b10000101 : out <= 8'd64;
      8'b11111010 : out <= 8'd65;
      8'b01111101 : out <= 8'd66;
      8'b10000110 : out <= 8'd67;
      8'b01000011 : out <= 8'd68;
      8'b10011001 : out <= 8'd69;
      8'b11110100 : out <= 8'd70;
      8'b01111010 : out <= 8'd71;
      8'b00111101 : out <= 8'd72;
      8'b10100110 : out <= 8'd73;
      8'b01010011 : out <= 8'd74;
      8'b10010001 : out <= 8'd75;
      8'b11110000 : out <= 8'd76;
      8'b01111000 : out <= 8'd77;
      8'b00111100 : out <= 8'd78;
      8'b00011110 : out <= 8'd79;
      8'b00001111 : out <= 8'd80;
      8'b10111111 : out <= 8'd81;
      8'b11100111 : out <= 8'd82;
      8'b11001011 : out <= 8'd83;
      8'b11011101 : out <= 8'd84;
      8'b11010110 : out <= 8'd85;
      8'b01101011 : out <= 8'd86;
      8'b10001101 : out <= 8'd87;
      8'b11111110 : out <= 8'd88;
      8'b01111111 : out <= 8'd89;
      8'b10000111 : out <= 8'd90;
      8'b11111011 : out <= 8'd91;
      8'b11000101 : out <= 8'd92;
      8'b11011010 : out <= 8'd93;
      8'b01101101 : out <= 8'd94;
      8'b10001110 : out <= 8'd95;
      8'b01000111 : out <= 8'd96;
      8'b10011011 : out <= 8'd97;
      8'b11110101 : out <= 8'd98;
      8'b11000010 : out <= 8'd99;
      8'b01100001 : out <= 8'd100;
      8'b10001000 : out <= 8'd101;
      8'b01000100 : out <= 8'd102;
      8'b00100010 : out <= 8'd103;
      8'b00010001 : out <= 8'd104;
      8'b10110000 : out <= 8'd105;
      8'b01011000 : out <= 8'd106;
      8'b00101100 : out <= 8'd107;
      8'b00010110 : out <= 8'd108;
      8'b00001011 : out <= 8'd109;
      8'b10111101 : out <= 8'd110;
      8'b11100110 : out <= 8'd111;
      8'b01110011 : out <= 8'd112;
      8'b10000001 : out <= 8'd113;
      8'b11111000 : out <= 8'd114;
      8'b01111100 : out <= 8'd115;
      8'b00111110 : out <= 8'd116;
      8'b00011111 : out <= 8'd117;
      8'b10110111 : out <= 8'd118;
      8'b11100011 : out <= 8'd119;
      8'b11001001 : out <= 8'd120;
      8'b11011100 : out <= 8'd121;
      8'b01101110 : out <= 8'd122;
      8'b00110111 : out <= 8'd123;
      8'b10100011 : out <= 8'd124;
      8'b11101001 : out <= 8'd125;
      8'b11001100 : out <= 8'd126;
      8'b01100110 : out <= 8'd127;
      8'b00110011 : out <= 8'd128;
      8'b10100001 : out <= 8'd129;
      8'b11101000 : out <= 8'd130;
      8'b01110100 : out <= 8'd131;
      8'b00111010 : out <= 8'd132;
      8'b00011101 : out <= 8'd133;
      8'b10110110 : out <= 8'd134;
      8'b01011011 : out <= 8'd135;
      8'b10010101 : out <= 8'd136;
      8'b11110010 : out <= 8'd137;
      8'b01111001 : out <= 8'd138;
      8'b10000100 : out <= 8'd139;
      8'b01000010 : out <= 8'd140;
      8'b00100001 : out <= 8'd141;
      8'b10101000 : out <= 8'd142;
      8'b01010100 : out <= 8'd143;
      8'b00101010 : out <= 8'd144;
      8'b00010101 : out <= 8'd145;
      8'b10110010 : out <= 8'd146;
      8'b01011001 : out <= 8'd147;
      8'b10010100 : out <= 8'd148;
      8'b01001010 : out <= 8'd149;
      8'b00100101 : out <= 8'd150;
      8'b10101010 : out <= 8'd151;
      8'b01010101 : out <= 8'd152;
      8'b10010010 : out <= 8'd153;
      8'b01001001 : out <= 8'd154;
      8'b10011100 : out <= 8'd155;
      8'b01001110 : out <= 8'd156;
      8'b00100111 : out <= 8'd157;
      8'b10101011 : out <= 8'd158;
      8'b11101101 : out <= 8'd159;
      8'b11001110 : out <= 8'd160;
      8'b01100111 : out <= 8'd161;
      8'b10001011 : out <= 8'd162;
      8'b11111101 : out <= 8'd163;
      8'b11000110 : out <= 8'd164;
      8'b01100011 : out <= 8'd165;
      8'b10001001 : out <= 8'd166;
      8'b11111100 : out <= 8'd167;
      8'b01111110 : out <= 8'd168;
      8'b00111111 : out <= 8'd169;
      8'b10100111 : out <= 8'd170;
      8'b11101011 : out <= 8'd171;
      8'b11001101 : out <= 8'd172;
      8'b11011110 : out <= 8'd173;
      8'b01101111 : out <= 8'd174;
      8'b10001111 : out <= 8'd175;
      8'b11111111 : out <= 8'd176;
      8'b11000111 : out <= 8'd177;
      8'b11011011 : out <= 8'd178;
      8'b11010101 : out <= 8'd179;
      8'b11010010 : out <= 8'd180;
      8'b01101001 : out <= 8'd181;
      8'b10001100 : out <= 8'd182;
      8'b01000110 : out <= 8'd183;
      8'b00100011 : out <= 8'd184;
      8'b10101001 : out <= 8'd185;
      8'b11101100 : out <= 8'd186;
      8'b01110110 : out <= 8'd187;
      8'b00111011 : out <= 8'd188;
      8'b10100101 : out <= 8'd189;
      8'b11101010 : out <= 8'd190;
      8'b01110101 : out <= 8'd191;
      8'b10000010 : out <= 8'd192;
      8'b01000001 : out <= 8'd193;
      8'b10011000 : out <= 8'd194;
      8'b01001100 : out <= 8'd195;
      8'b00100110 : out <= 8'd196;
      8'b00010011 : out <= 8'd197;
      8'b10110001 : out <= 8'd198;
      8'b11100000 : out <= 8'd199;
      8'b01110000 : out <= 8'd200;
      8'b00111000 : out <= 8'd201;
      8'b00011100 : out <= 8'd202;
      8'b00001110 : out <= 8'd203;
      8'b00000111 : out <= 8'd204;
      8'b10111011 : out <= 8'd205;
      8'b11100101 : out <= 8'd206;
      8'b11001010 : out <= 8'd207;
      8'b01100101 : out <= 8'd208;
      8'b10001010 : out <= 8'd209;
      8'b01000101 : out <= 8'd210;
      8'b10011010 : out <= 8'd211;
      8'b01001101 : out <= 8'd212;
      8'b10011110 : out <= 8'd213;
      8'b01001111 : out <= 8'd214;
      8'b10011111 : out <= 8'd215;
      8'b11110111 : out <= 8'd216;
      8'b11000011 : out <= 8'd217;
      8'b11011001 : out <= 8'd218;
      8'b11010100 : out <= 8'd219;
      8'b01101010 : out <= 8'd220;
      8'b00110101 : out <= 8'd221;
      8'b10100010 : out <= 8'd222;
      8'b01010001 : out <= 8'd223;
      8'b10010000 : out <= 8'd224;
      8'b01001000 : out <= 8'd225;
      8'b00100100 : out <= 8'd226;
      8'b00010010 : out <= 8'd227;
      8'b00001001 : out <= 8'd228;
      8'b10111100 : out <= 8'd229;
      8'b01011110 : out <= 8'd230;
      8'b00101111 : out <= 8'd231;
      8'b10101111 : out <= 8'd232;
      8'b11101111 : out <= 8'd233;
      8'b11001111 : out <= 8'd234;
      8'b11011111 : out <= 8'd235;
      8'b11010111 : out <= 8'd236;
      8'b11010011 : out <= 8'd237;
      8'b11010001 : out <= 8'd238;
      8'b11010000 : out <= 8'd239;
      8'b01101000 : out <= 8'd240;
      8'b00110100 : out <= 8'd241;
      8'b00011010 : out <= 8'd242;
      8'b00001101 : out <= 8'd243;
      8'b10111110 : out <= 8'd244;
      8'b01011111 : out <= 8'd245;
      8'b10010111 : out <= 8'd246;
      8'b11110011 : out <= 8'd247;
      8'b11000001 : out <= 8'd248;
      8'b11011000 : out <= 8'd249;
      8'b01101100 : out <= 8'd250;
      8'b00110110 : out <= 8'd251;
      8'b00011011 : out <= 8'd252;
      8'b10110101 : out <= 8'd253;
      8'b11100010 : out <= 8'd254;
      8'b01110001 : out <= 8'd255;
      default: out <= 8'd0;
    endcase
  end
endmodule

