`define SYMBOL_WIDTH 8
`define N 18
`define K 16


module RS_Encoder
(
  input wire [(`SYMBOL_WIDTH * `K)-1:0] in,
  output wire [(`SYMBOL_WIDTH * `N)-1:0] out
);
  
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_0;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_1;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_2;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_3;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_4;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_5;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_6;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_7;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_8;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_9;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_10;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_11;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_12;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_13;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_14;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_15;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_16;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_17;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_18;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_19;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_20;
  wire  [(`SYMBOL_WIDTH * `N):0] G_row_21;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_22;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_23;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_24;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_25;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_26;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_27;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_28;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_29;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_30;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_31;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_32;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_33;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_34;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_35;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_36;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_37;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_38;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_39;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_40;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_41;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_42;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_43;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_44;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_45;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_46;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_47;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_48;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_49;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_50;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_51;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_52;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_53;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_54;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_55;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_56;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_57;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_58;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_59;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_60;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_61;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_62;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_63;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_64;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_65;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_66;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_67;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_68;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_69;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_70;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_71;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_72;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_73;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_74;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_75;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_76;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_77;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_78;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_79;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_80;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_81;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_82;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_83;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_84;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_85;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_86;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_87;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_88;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_89;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_90;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_91;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_92;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_93;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_94;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_95;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_96;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_97;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_98;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_99;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_100;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_101;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_102;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_103;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_104;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_105;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_106;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_107;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_108;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_109;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_110;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_111;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_112;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_113;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_114;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_115;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_116;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_117;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_118;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_119;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_120;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_121;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_122;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_123;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_124;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_125;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_126;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_127;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_128;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_129;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_130;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_131;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_132;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_133;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_134;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_135;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_136;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_137;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_138;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_139;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_140;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_141;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_142;
wire  [(`SYMBOL_WIDTH * `N):0] G_row_143;

  
assign G_row_0 = 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_1 = 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_2 = 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_3 = 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_4 = 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_5 = 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_6 = 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_7 = 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_8 = 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_9 = 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_10 = 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_11 = 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_12 = 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_13 = 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_14 = 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_15 = 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_16 = 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_17 = 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_18 = 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_19 = 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_20 = 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_21 = 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_22 = 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_23 = 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_24 = 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_25 = 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_26 = 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_27 = 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_28 = 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_29 = 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_30 = 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_31 = 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_32 = 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_33 = 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_34 = 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_35 = 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_36 = 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_37 = 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_38 = 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_39 = 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_40 = 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_41 = 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_42 = 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_43 = 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_44 = 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_45 = 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_46 = 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_47 = 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_48 = 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_49 = 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_50 = 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_51 = 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_52 = 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_53 = 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_54 = 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_55 = 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_56 = 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_57 = 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_58 = 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_59 = 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_60 = 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_61 = 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
assign G_row_62 = 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
assign G_row_63 = 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
assign G_row_64 = 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
assign G_row_65 = 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
assign G_row_66 = 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
assign G_row_67 = 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
assign G_row_68 = 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
assign G_row_69 = 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
assign G_row_70 = 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
assign G_row_71 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
assign G_row_72 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
assign G_row_73 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
assign G_row_74 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
assign G_row_75 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
assign G_row_76 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
assign G_row_77 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
assign G_row_78 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
assign G_row_79 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
assign G_row_80 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
assign G_row_81 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
assign G_row_82 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
assign G_row_83 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
assign G_row_84 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
assign G_row_85 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
assign G_row_86 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
assign G_row_87 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
assign G_row_88 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
assign G_row_89 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
assign G_row_90 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
assign G_row_91 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
assign G_row_92 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
assign G_row_93 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
assign G_row_94 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
assign G_row_95 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
assign G_row_96 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
assign G_row_97 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
assign G_row_98 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
assign G_row_99 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
assign G_row_100 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
assign G_row_101 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
assign G_row_102 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
assign G_row_103 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
assign G_row_104 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
assign G_row_105 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
assign G_row_106 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
assign G_row_107 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
assign G_row_108 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
assign G_row_109 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
assign G_row_110 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
assign G_row_111 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
assign G_row_112 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
assign G_row_113 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
assign G_row_114 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
assign G_row_115 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
assign G_row_116 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
assign G_row_117 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
assign G_row_118 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
assign G_row_119 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
assign G_row_120 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
assign G_row_121 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
assign G_row_122 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
assign G_row_123 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
assign G_row_124 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
assign G_row_125 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
assign G_row_126 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
assign G_row_127 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
assign G_row_128 = 128'b01000111111010111000011110111111101000000110111110111000000111111101111110011011111100000111011111011000001101000000110000000011;
assign G_row_129 = 128'b00100011011101010100001101011111010100001011011101011100000011110110111111001101111110001011101101101100000110100000011010000001;
assign G_row_130 = 128'b10010001101110101010000100101111101010001101101110101110100001111011011111100110011111001101110100110110000011011000001111000000;
assign G_row_131 = 128'b01001000010111011101000010010111110101001110110101010111010000111101101111110011101111100110111000011011100001101100000101100000;
assign G_row_132 = 128'b11100011110001010110111101110100110010101001100100010011101111100011001011100010001011110100000001010101111101111110110000110011;
assign G_row_133 = 128'b10110110100010010011000010000101010001011010001110110001110000000100011011101010011001110101011101110010110011110111101000011010;
assign G_row_134 = 128'b00011100101011110001111111111101100000101011111011100000011111110111110001101110110000111101110001100001110100110011000100001110;
assign G_row_135 = 128'b10001110110101110000111101111110010000011101111101110000001111111011111000110111111000011110111010110000011010010001100000000111;
assign G_row_136 = 128'b01011110001111111111101100000100011111001100000111111111111110001101110110000110101110011100001010100110011000100001110100000101;
assign G_row_137 = 128'b10101111000111111111110110000010101111101110000001111111011111000110111011000011110111000110000111010011001100010000111000000010;
assign G_row_138 = 128'b11010111000011110111111001000001110111110111000000111111101111100011011111100001111011101011000001101001000110000000011100000001;
assign G_row_139 = 128'b11101011100001111011111110100000011011111011100000011111110111111001101111110000011101111101100000110100000011000000001110000000;
assign G_row_140 = 128'b00101011011111001010010001010100110010111001110111110000100101110001000001111110000000101010111010111100011001001001110001000101;
assign G_row_141 = 128'b01001011100000010010100100101110000110011000111100000111001100110101010100111001101110001001010101111000110100001101001100100111;
assign G_row_142 = 128'b01111011111111111110111100010011111100000000011011111100111000010111011100011010111001010000100010011010100010100111010000010110;
assign G_row_143 = 128'b10111101011111111111011100001001111110001000001111111110111100001011101100001101011100101000010001001101110001010011101000001011;
  
assign out[143]  =^(in & G_row_0) ;
assign out[142]  =^(in & G_row_1) ;
assign out[141]  =^(in & G_row_2) ;
assign out[140]  =^(in & G_row_3) ;
assign out[139]  =^(in & G_row_4) ;
assign out[138]  =^(in & G_row_5) ;
assign out[137]  =^(in & G_row_6) ;
assign out[136]  =^(in & G_row_7) ;
assign out[135]  =^(in & G_row_8) ;
assign out[134]  =^(in & G_row_9) ;
assign out[133]  =^(in & G_row_10) ;
assign out[132]  =^(in & G_row_11) ;
assign out[131]  =^(in & G_row_12) ;
assign out[130]  =^(in & G_row_13) ;
assign out[129]  =^(in & G_row_14) ;
assign out[128]  =^(in & G_row_15) ;
assign out[127]  =^(in & G_row_16) ;
assign out[126]  =^(in & G_row_17) ;
assign out[125]  =^(in & G_row_18) ;
assign out[124]  =^(in & G_row_19) ;
assign out[123]  =^(in & G_row_20) ;
assign out[122]  =^(in & G_row_21) ;
assign out[121]  =^(in & G_row_22) ;
assign out[120]  =^(in & G_row_23) ;
assign out[119]  =^(in & G_row_24) ;
assign out[118]  =^(in & G_row_25) ;
assign out[117]  =^(in & G_row_26) ;
assign out[116]  =^(in & G_row_27) ;
assign out[115]  =^(in & G_row_28) ;
assign out[114]  =^(in & G_row_29) ;
assign out[113]  =^(in & G_row_30) ;
assign out[112]  =^(in & G_row_31) ;
assign out[111]  =^(in & G_row_32) ;
assign out[110]  =^(in & G_row_33) ;
assign out[109]  =^(in & G_row_34) ;
assign out[108]  =^(in & G_row_35) ;
assign out[107]  =^(in & G_row_36) ;
assign out[106]  =^(in & G_row_37) ;
assign out[105]  =^(in & G_row_38) ;
assign out[104]  =^(in & G_row_39) ;
assign out[103]  =^(in & G_row_40) ;
assign out[102]  =^(in & G_row_41) ;
assign out[101]  =^(in & G_row_42) ;
assign out[100]  =^(in & G_row_43) ;
assign out[99]  =^(in & G_row_44) ;
assign out[98]  =^(in & G_row_45) ;
assign out[97]  =^(in & G_row_46) ;
assign out[96]  =^(in & G_row_47) ;
assign out[95]  =^(in & G_row_48) ;
assign out[94]  =^(in & G_row_49) ;
assign out[93]  =^(in & G_row_50) ;
assign out[92]  =^(in & G_row_51) ;
assign out[91]  =^(in & G_row_52) ;
assign out[90]  =^(in & G_row_53) ;
assign out[89]  =^(in & G_row_54) ;
assign out[88]  =^(in & G_row_55) ;
assign out[87]  =^(in & G_row_56) ;
assign out[86]  =^(in & G_row_57) ;
assign out[85]  =^(in & G_row_58) ;
assign out[84]  =^(in & G_row_59) ;
assign out[83]  =^(in & G_row_60) ;
assign out[82]  =^(in & G_row_61) ;
assign out[81]  =^(in & G_row_62) ;
assign out[80]  =^(in & G_row_63) ;
assign out[79]  =^(in & G_row_64) ;
assign out[78]  =^(in & G_row_65) ;
assign out[77]  =^(in & G_row_66) ;
assign out[76]  =^(in & G_row_67) ;
assign out[75]  =^(in & G_row_68) ;
assign out[74]  =^(in & G_row_69) ;
assign out[73]  =^(in & G_row_70) ;
assign out[72]  =^(in & G_row_71) ;
assign out[71]  =^(in & G_row_72) ;
assign out[70]  =^(in & G_row_73) ;
assign out[69]  =^(in & G_row_74) ;
assign out[68]  =^(in & G_row_75) ;
assign out[67]  =^(in & G_row_76) ;
assign out[66]  =^(in & G_row_77) ;
assign out[65]  =^(in & G_row_78) ;
assign out[64]  =^(in & G_row_79) ;
assign out[63]  =^(in & G_row_80) ;
assign out[62]  =^(in & G_row_81) ;
assign out[61]  =^(in & G_row_82) ;
assign out[60]  =^(in & G_row_83) ;
assign out[59]  =^(in & G_row_84) ;
assign out[58]  =^(in & G_row_85) ;
assign out[57]  =^(in & G_row_86) ;
assign out[56]  =^(in & G_row_87) ;
assign out[55]  =^(in & G_row_88) ;
assign out[54]  =^(in & G_row_89) ;
assign out[53]  =^(in & G_row_90) ;
assign out[52]  =^(in & G_row_91) ;
assign out[51]  =^(in & G_row_92) ;
assign out[50]  =^(in & G_row_93) ;
assign out[49]  =^(in & G_row_94) ;
assign out[48]  =^(in & G_row_95) ;
assign out[47]  =^(in & G_row_96) ;
assign out[46]  =^(in & G_row_97) ;
assign out[45]  =^(in & G_row_98) ;
assign out[44]  =^(in & G_row_99) ;
assign out[43]  =^(in & G_row_100) ;
assign out[42]  =^(in & G_row_101) ;
assign out[41]  =^(in & G_row_102) ;
assign out[40]  =^(in & G_row_103) ;
assign out[39]  =^(in & G_row_104) ;
assign out[38]  =^(in & G_row_105) ;
assign out[37]  =^(in & G_row_106) ;
assign out[36]  =^(in & G_row_107) ;
assign out[35]  =^(in & G_row_108) ;
assign out[34]  =^(in & G_row_109) ;
assign out[33]  =^(in & G_row_110) ;
assign out[32]  =^(in & G_row_111) ;
assign out[31]  =^(in & G_row_112) ;
assign out[30]  =^(in & G_row_113) ;
assign out[29]  =^(in & G_row_114) ;
assign out[28]  =^(in & G_row_115) ;
assign out[27]  =^(in & G_row_116) ;
assign out[26]  =^(in & G_row_117) ;
assign out[25]  =^(in & G_row_118) ;
assign out[24]  =^(in & G_row_119) ;
assign out[23]  =^(in & G_row_120) ;
assign out[22]  =^(in & G_row_121) ;
assign out[21]  =^(in & G_row_122) ;
assign out[20]  =^(in & G_row_123) ;
assign out[19]  =^(in & G_row_124) ;
assign out[18]  =^(in & G_row_125) ;
assign out[17]  =^(in & G_row_126) ;
assign out[16]  =^(in & G_row_127) ;
assign out[15]  =^(in & G_row_128) ;
assign out[14]  =^(in & G_row_129) ;
assign out[13]  =^(in & G_row_130) ;
assign out[12]  =^(in & G_row_131) ;
assign out[11]  =^(in & G_row_132) ;
assign out[10]  =^(in & G_row_133) ;
assign out[9]  =^(in & G_row_134) ;
assign out[8]  =^(in & G_row_135) ;
assign out[7]  =^(in & G_row_136) ;
assign out[6]  =^(in & G_row_137) ;
assign out[5]  =^(in & G_row_138) ;
assign out[4]  =^(in & G_row_139) ;
assign out[3]  =^(in & G_row_140) ;
assign out[2]  =^(in & G_row_141) ;
assign out[1]  =^(in & G_row_142) ;
assign out[0]  =^(in & G_row_143) ;
  
  
endmodule

