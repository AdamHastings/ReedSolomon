function bit [`SYMBOL_WIDTH-1:0] getSymbol (input int a);
  bit [`SYMBOL_WIDTH-1:0] s;

      if (a == 0) begin s=8'b00000000; end
      else if (a == 1) begin s=8'b10000000; end
      else if (a == 2) begin s=8'b01000000; end
      else if (a == 3) begin s=8'b00100000; end
      else if (a == 4) begin s=8'b00010000; end
      else if (a == 5) begin s=8'b00001000; end
      else if (a == 6) begin s=8'b00000100; end
      else if (a == 7) begin s=8'b00000010; end
      else if (a == 8) begin s=8'b00000001; end
      else if (a == 9) begin s=8'b10111000; end
      else if (a == 10) begin s=8'b01011100; end
      else if (a == 11) begin s=8'b00101110; end
      else if (a == 12) begin s=8'b00010111; end
      else if (a == 13) begin s=8'b10110011; end
      else if (a == 14) begin s=8'b11100001; end
      else if (a == 15) begin s=8'b11001000; end
      else if (a == 16) begin s=8'b01100100; end
      else if (a == 17) begin s=8'b00110010; end
      else if (a == 18) begin s=8'b00011001; end
      else if (a == 19) begin s=8'b10110100; end
      else if (a == 20) begin s=8'b01011010; end
      else if (a == 21) begin s=8'b00101101; end
      else if (a == 22) begin s=8'b10101110; end
      else if (a == 23) begin s=8'b01010111; end
      else if (a == 24) begin s=8'b10010011; end
      else if (a == 25) begin s=8'b11110001; end
      else if (a == 26) begin s=8'b11000000; end
      else if (a == 27) begin s=8'b01100000; end
      else if (a == 28) begin s=8'b00110000; end
      else if (a == 29) begin s=8'b00011000; end
      else if (a == 30) begin s=8'b00001100; end
      else if (a == 31) begin s=8'b00000110; end
      else if (a == 32) begin s=8'b00000011; end
      else if (a == 33) begin s=8'b10111001; end
      else if (a == 34) begin s=8'b11100100; end
      else if (a == 35) begin s=8'b01110010; end
      else if (a == 36) begin s=8'b00111001; end
      else if (a == 37) begin s=8'b10100100; end
      else if (a == 38) begin s=8'b01010010; end
      else if (a == 39) begin s=8'b00101001; end
      else if (a == 40) begin s=8'b10101100; end
      else if (a == 41) begin s=8'b01010110; end
      else if (a == 42) begin s=8'b00101011; end
      else if (a == 43) begin s=8'b10101101; end
      else if (a == 44) begin s=8'b11101110; end
      else if (a == 45) begin s=8'b01110111; end
      else if (a == 46) begin s=8'b10000011; end
      else if (a == 47) begin s=8'b11111001; end
      else if (a == 48) begin s=8'b11000100; end
      else if (a == 49) begin s=8'b01100010; end
      else if (a == 50) begin s=8'b00110001; end
      else if (a == 51) begin s=8'b10100000; end
      else if (a == 52) begin s=8'b01010000; end
      else if (a == 53) begin s=8'b00101000; end
      else if (a == 54) begin s=8'b00010100; end
      else if (a == 55) begin s=8'b00001010; end
      else if (a == 56) begin s=8'b00000101; end
      else if (a == 57) begin s=8'b10111010; end
      else if (a == 58) begin s=8'b01011101; end
      else if (a == 59) begin s=8'b10010110; end
      else if (a == 60) begin s=8'b01001011; end
      else if (a == 61) begin s=8'b10011101; end
      else if (a == 62) begin s=8'b11110110; end
      else if (a == 63) begin s=8'b01111011; end
      else if (a == 64) begin s=8'b10000101; end
      else if (a == 65) begin s=8'b11111010; end
      else if (a == 66) begin s=8'b01111101; end
      else if (a == 67) begin s=8'b10000110; end
      else if (a == 68) begin s=8'b01000011; end
      else if (a == 69) begin s=8'b10011001; end
      else if (a == 70) begin s=8'b11110100; end
      else if (a == 71) begin s=8'b01111010; end
      else if (a == 72) begin s=8'b00111101; end
      else if (a == 73) begin s=8'b10100110; end
      else if (a == 74) begin s=8'b01010011; end
      else if (a == 75) begin s=8'b10010001; end
      else if (a == 76) begin s=8'b11110000; end
      else if (a == 77) begin s=8'b01111000; end
      else if (a == 78) begin s=8'b00111100; end
      else if (a == 79) begin s=8'b00011110; end
      else if (a == 80) begin s=8'b00001111; end
      else if (a == 81) begin s=8'b10111111; end
      else if (a == 82) begin s=8'b11100111; end
      else if (a == 83) begin s=8'b11001011; end
      else if (a == 84) begin s=8'b11011101; end
      else if (a == 85) begin s=8'b11010110; end
      else if (a == 86) begin s=8'b01101011; end
      else if (a == 87) begin s=8'b10001101; end
      else if (a == 88) begin s=8'b11111110; end
      else if (a == 89) begin s=8'b01111111; end
      else if (a == 90) begin s=8'b10000111; end
      else if (a == 91) begin s=8'b11111011; end
      else if (a == 92) begin s=8'b11000101; end
      else if (a == 93) begin s=8'b11011010; end
      else if (a == 94) begin s=8'b01101101; end
      else if (a == 95) begin s=8'b10001110; end
      else if (a == 96) begin s=8'b01000111; end
      else if (a == 97) begin s=8'b10011011; end
      else if (a == 98) begin s=8'b11110101; end
      else if (a == 99) begin s=8'b11000010; end
      else if (a == 100) begin s=8'b01100001; end
      else if (a == 101) begin s=8'b10001000; end
      else if (a == 102) begin s=8'b01000100; end
      else if (a == 103) begin s=8'b00100010; end
      else if (a == 104) begin s=8'b00010001; end
      else if (a == 105) begin s=8'b10110000; end
      else if (a == 106) begin s=8'b01011000; end
      else if (a == 107) begin s=8'b00101100; end
      else if (a == 108) begin s=8'b00010110; end
      else if (a == 109) begin s=8'b00001011; end
      else if (a == 110) begin s=8'b10111101; end
      else if (a == 111) begin s=8'b11100110; end
      else if (a == 112) begin s=8'b01110011; end
      else if (a == 113) begin s=8'b10000001; end
      else if (a == 114) begin s=8'b11111000; end
      else if (a == 115) begin s=8'b01111100; end
      else if (a == 116) begin s=8'b00111110; end
      else if (a == 117) begin s=8'b00011111; end
      else if (a == 118) begin s=8'b10110111; end
      else if (a == 119) begin s=8'b11100011; end
      else if (a == 120) begin s=8'b11001001; end
      else if (a == 121) begin s=8'b11011100; end
      else if (a == 122) begin s=8'b01101110; end
      else if (a == 123) begin s=8'b00110111; end
      else if (a == 124) begin s=8'b10100011; end
      else if (a == 125) begin s=8'b11101001; end
      else if (a == 126) begin s=8'b11001100; end
      else if (a == 127) begin s=8'b01100110; end
      else if (a == 128) begin s=8'b00110011; end
      else if (a == 129) begin s=8'b10100001; end
      else if (a == 130) begin s=8'b11101000; end
      else if (a == 131) begin s=8'b01110100; end
      else if (a == 132) begin s=8'b00111010; end
      else if (a == 133) begin s=8'b00011101; end
      else if (a == 134) begin s=8'b10110110; end
      else if (a == 135) begin s=8'b01011011; end
      else if (a == 136) begin s=8'b10010101; end
      else if (a == 137) begin s=8'b11110010; end
      else if (a == 138) begin s=8'b01111001; end
      else if (a == 139) begin s=8'b10000100; end
      else if (a == 140) begin s=8'b01000010; end
      else if (a == 141) begin s=8'b00100001; end
      else if (a == 142) begin s=8'b10101000; end
      else if (a == 143) begin s=8'b01010100; end
      else if (a == 144) begin s=8'b00101010; end
      else if (a == 145) begin s=8'b00010101; end
      else if (a == 146) begin s=8'b10110010; end
      else if (a == 147) begin s=8'b01011001; end
      else if (a == 148) begin s=8'b10010100; end
      else if (a == 149) begin s=8'b01001010; end
      else if (a == 150) begin s=8'b00100101; end
      else if (a == 151) begin s=8'b10101010; end
      else if (a == 152) begin s=8'b01010101; end
      else if (a == 153) begin s=8'b10010010; end
      else if (a == 154) begin s=8'b01001001; end
      else if (a == 155) begin s=8'b10011100; end
      else if (a == 156) begin s=8'b01001110; end
      else if (a == 157) begin s=8'b00100111; end
      else if (a == 158) begin s=8'b10101011; end
      else if (a == 159) begin s=8'b11101101; end
      else if (a == 160) begin s=8'b11001110; end
      else if (a == 161) begin s=8'b01100111; end
      else if (a == 162) begin s=8'b10001011; end
      else if (a == 163) begin s=8'b11111101; end
      else if (a == 164) begin s=8'b11000110; end
      else if (a == 165) begin s=8'b01100011; end
      else if (a == 166) begin s=8'b10001001; end
      else if (a == 167) begin s=8'b11111100; end
      else if (a == 168) begin s=8'b01111110; end
      else if (a == 169) begin s=8'b00111111; end
      else if (a == 170) begin s=8'b10100111; end
      else if (a == 171) begin s=8'b11101011; end
      else if (a == 172) begin s=8'b11001101; end
      else if (a == 173) begin s=8'b11011110; end
      else if (a == 174) begin s=8'b01101111; end
      else if (a == 175) begin s=8'b10001111; end
      else if (a == 176) begin s=8'b11111111; end
      else if (a == 177) begin s=8'b11000111; end
      else if (a == 178) begin s=8'b11011011; end
      else if (a == 179) begin s=8'b11010101; end
      else if (a == 180) begin s=8'b11010010; end
      else if (a == 181) begin s=8'b01101001; end
      else if (a == 182) begin s=8'b10001100; end
      else if (a == 183) begin s=8'b01000110; end
      else if (a == 184) begin s=8'b00100011; end
      else if (a == 185) begin s=8'b10101001; end
      else if (a == 186) begin s=8'b11101100; end
      else if (a == 187) begin s=8'b01110110; end
      else if (a == 188) begin s=8'b00111011; end
      else if (a == 189) begin s=8'b10100101; end
      else if (a == 190) begin s=8'b11101010; end
      else if (a == 191) begin s=8'b01110101; end
      else if (a == 192) begin s=8'b10000010; end
      else if (a == 193) begin s=8'b01000001; end
      else if (a == 194) begin s=8'b10011000; end
      else if (a == 195) begin s=8'b01001100; end
      else if (a == 196) begin s=8'b00100110; end
      else if (a == 197) begin s=8'b00010011; end
      else if (a == 198) begin s=8'b10110001; end
      else if (a == 199) begin s=8'b11100000; end
      else if (a == 200) begin s=8'b01110000; end
      else if (a == 201) begin s=8'b00111000; end
      else if (a == 202) begin s=8'b00011100; end
      else if (a == 203) begin s=8'b00001110; end
      else if (a == 204) begin s=8'b00000111; end
      else if (a == 205) begin s=8'b10111011; end
      else if (a == 206) begin s=8'b11100101; end
      else if (a == 207) begin s=8'b11001010; end
      else if (a == 208) begin s=8'b01100101; end
      else if (a == 209) begin s=8'b10001010; end
      else if (a == 210) begin s=8'b01000101; end
      else if (a == 211) begin s=8'b10011010; end
      else if (a == 212) begin s=8'b01001101; end
      else if (a == 213) begin s=8'b10011110; end
      else if (a == 214) begin s=8'b01001111; end
      else if (a == 215) begin s=8'b10011111; end
      else if (a == 216) begin s=8'b11110111; end
      else if (a == 217) begin s=8'b11000011; end
      else if (a == 218) begin s=8'b11011001; end
      else if (a == 219) begin s=8'b11010100; end
      else if (a == 220) begin s=8'b01101010; end
      else if (a == 221) begin s=8'b00110101; end
      else if (a == 222) begin s=8'b10100010; end
      else if (a == 223) begin s=8'b01010001; end
      else if (a == 224) begin s=8'b10010000; end
      else if (a == 225) begin s=8'b01001000; end
      else if (a == 226) begin s=8'b00100100; end
      else if (a == 227) begin s=8'b00010010; end
      else if (a == 228) begin s=8'b00001001; end
      else if (a == 229) begin s=8'b10111100; end
      else if (a == 230) begin s=8'b01011110; end
      else if (a == 231) begin s=8'b00101111; end
      else if (a == 232) begin s=8'b10101111; end
      else if (a == 233) begin s=8'b11101111; end
      else if (a == 234) begin s=8'b11001111; end
      else if (a == 235) begin s=8'b11011111; end
      else if (a == 236) begin s=8'b11010111; end
      else if (a == 237) begin s=8'b11010011; end
      else if (a == 238) begin s=8'b11010001; end
      else if (a == 239) begin s=8'b11010000; end
      else if (a == 240) begin s=8'b01101000; end
      else if (a == 241) begin s=8'b00110100; end
      else if (a == 242) begin s=8'b00011010; end
      else if (a == 243) begin s=8'b00001101; end
      else if (a == 244) begin s=8'b10111110; end
      else if (a == 245) begin s=8'b01011111; end
      else if (a == 246) begin s=8'b10010111; end
      else if (a == 247) begin s=8'b11110011; end
      else if (a == 248) begin s=8'b11000001; end
      else if (a == 249) begin s=8'b11011000; end
      else if (a == 250) begin s=8'b01101100; end
      else if (a == 251) begin s=8'b00110110; end
      else if (a == 252) begin s=8'b00011011; end
      else if (a == 253) begin s=8'b10110101; end
      else if (a == 254) begin s=8'b11100010; end
      else if (a == 255) begin s=8'b01110001; end

      return s;
    
endfunction
